library verilog;
use verilog.vl_types.all;
entity procfixcba_tb is
end procfixcba_tb;
